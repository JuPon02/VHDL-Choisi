ibrary IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LED is
	port(
		 );
end entity;

architecture rtl of LED is
	begin
		
end rtl;