ibrary IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Switch is
	port(
	
		 );
end entity;

architecture rtl of Switch is
	begin
		
end rtl;