ibrary IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Random is
	port(
		 );
end entity;

architecture rtl of Random is
	begin
		
end rtl;
--test